-- =============================================================================
-- AUTHOR:          Le Vu Duc Hung
--
-- DATE:            13/06/2023
--
-- FILE:            adc_pkg.vhd
-- =============================================================================
-- MIT License
-- Copyright (c) 2023 Le Vu Duc Hung
--
-- Permission is hereby granted, free of charge, to any person obtaining
-- a copy of this software and associated documentation files (the
-- "Software"), to deal in the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
--
-- The above copyright notice and this permission notice shall be
-- included in all copies or substantial portions of the Software.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND,
-- EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND
-- NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS BE
-- LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION
-- OF CONTRACT, TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION
-- WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE SOFTWARE.
-- =============================================================================

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package adc_pkg is

    --================================= Types =====================================--
    type adc_config is record
        clock_frequency:        positive;  -- clock frequency (50MHz)
        data_bits:              positive;  -- Number of data bits per frame
        end_reception_state:    positive; 
        clk_div:                positive;
        ratio_must_be_half:     boolean;
        sampling_div:           positive;
    end record adc_config;
    

    --================================= Constants =================================--
    constant adc_default_config: adc_config := (
        clock_frequency         =>    50000000,
        data_bits               =>    8,
        end_reception_state     =>    12,
        clk_div                 =>    125,
        ratio_must_be_half      =>    false,
        sampling_div            =>    40
    );


    --===================================== ADC ====================================--
    component adc is
        
    end component adc;

end package adc_pkg;

package body adc_pkg is
       

end package body adc_pkg;
